module packet_dut;
endmodule
